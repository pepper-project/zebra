../../common/rtl/field_one_minus.sv