../../common/tb/prover_layer_test.sv