../../common/rtl/prover_compute_v.sv