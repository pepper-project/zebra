../../common/tb/prover_compute_v_test.sv