../../common/tb/simple_adder_tree_test.sv