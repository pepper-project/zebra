../../common/rtl/pergate_compute.sv