../../common/tb/prover_compute_h_test.sv