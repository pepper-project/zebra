../../common/rtl/field_arith_ns.sv