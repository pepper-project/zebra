../../common/rtl/prover_layer.sv