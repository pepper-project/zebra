../../common/tb/layer_declaration_test.sv