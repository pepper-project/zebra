../../common/rtl/verifier_interface_w0.sv