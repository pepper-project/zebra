../../common/rtl/verifier_interface.sv