../../common/tb/prover_verifier_test.sv