../../common/rtl/pergate_compute_fj.sv