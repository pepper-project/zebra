../../common/rtl/pergate_compute_seq.sv