../../common/rtl/computation_gatefn.sv