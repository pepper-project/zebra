../../common/rtl/computation_layer.sv