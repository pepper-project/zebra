../../common/tb/pergate_compute_test.sv