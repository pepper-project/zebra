../../common/rtl/prover_compute_h_elem.sv