../../common/rtl/prover_compute_w0_elem.sv