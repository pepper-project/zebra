../../common/rtl/prover_compute_w0.sv