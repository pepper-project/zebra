../../common/rtl/field_negate_or_double.sv