../../common/rtl/field_negate.sv