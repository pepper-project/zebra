../../common/tb/cmt_top_test.sv