../../common/rtl/layer_top.sv