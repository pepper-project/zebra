../../common/rtl/layer_top_pl.sv