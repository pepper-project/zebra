../../common/rtl/prover_compute_v_elem.sv