../../common/tb/field_arith_test.sv