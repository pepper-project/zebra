../../common/rtl/layer_ringbuf_pl.sv