../../common/tb/sram_generic_test.sv