../../common/tb/prover_synth_test_tb.sv