../../common/rtl/sram_generic.sv