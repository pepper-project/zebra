../../common/rtl/prover_adder_tree_pl.sv