../../common/rtl/pergate_compute_addmul.sv