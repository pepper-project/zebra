../../common/rtl/field_mux.sv