../../common/rtl/prover_shuffle_v_elem.sv