../../common/rtl/pergate_compute_am_fj.sv