// hello.v
// testbench for hello VPI module
// (C) 2015 Riad S. Wahby <rsw@cs.nyu.edu>

`include "simulator.v"

module main;
    initial $hello;
endmodule
