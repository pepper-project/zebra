../../common/rtl/prover_shuffle_v.sv