../../common/rtl/field_double.sv