../../common/rtl/pergate_compute_gatefn.sv