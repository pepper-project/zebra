../../common/rtl/shiftreg_simple.sv