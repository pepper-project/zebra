../../common/rtl/field_multiplier.sv