../../common/rtl/field_adder.sv