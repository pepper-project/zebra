../../common/rtl/field_subtract.sv