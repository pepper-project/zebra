../../common/rtl/ringbuf_simple.sv