../../common/rtl/prover_compute_c012_fm1.sv