../../common/tb/prover_adder_tree_pl_test.sv