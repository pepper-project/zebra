../../common/tb/cmt_top_pl_test.sv