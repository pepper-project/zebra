../../common/rtl/prover_compute_h.sv