../../common/tb/prover_shuffle_v_test.sv