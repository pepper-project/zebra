../../common/rtl/pergate_compute_am012.sv