../../common/rtl/pergate_compute_gatefn_seq.sv